//A header file containing all the coefficients for the final product.

//for c1_scaled
localparam signed [55:0] C1_0  =  56'sd889574400;
localparam signed [55:0] C1_1  =  56'sd4670265600;
localparam signed [55:0] C1_2  = -56'sd6227020800;
localparam signed [55:0] C1_3  = -56'sd1297296000;
localparam signed [55:0] C1_4  =  56'sd2335132800;
localparam signed [55:0] C1_5  =  56'sd345945600;
localparam signed [55:0] C1_6  = -56'sd864864000;
localparam signed [55:0] C1_7  = -56'sd70761600;
localparam signed [55:0] C1_8  =  56'sd259459200;
localparam signed [55:0] C1_9  =  56'sd9434880;
localparam signed [55:0] C1_10 = -56'sd56609280;
localparam signed [55:0] C1_11 = -56'sd604800;
localparam signed [55:0] C1_12 =  56'sd7862400;
localparam signed [55:0] C1_13 = -56'sd518400;
localparam signed [55:0] C1_14 =  56'sd22596613079040000;

//for c2_scaled
localparam signed [52:0] C2_0  = -53'sd9286909632;
localparam signed [52:0] C2_1  =  53'sd5337446400;
localparam signed [52:0] C2_2  =  53'sd5337446400;
localparam signed [52:0] C2_3  = -53'sd833976000;
localparam signed [52:0] C2_4  = -53'sd833976000;
localparam signed [52:0] C2_5  =  53'sd164736000;
localparam signed [52:0] C2_6  =  53'sd164736000;
localparam signed [52:0] C2_7  = -53'sd27799200;
localparam signed [52:0] C2_8  = -53'sd27799200;
localparam signed [52:0] C2_9  =  53'sd3234816;
localparam signed [52:0] C2_10 =  53'sd3234816;
localparam signed [52:0] C2_11 = -53'sd187200;
localparam signed [52:0] C2_12 = -53'sd187200;
localparam signed [52:0] C2_14 =  53'sd3228087582720000;

//for c3_scaled
localparam signed [55:0] C3_0  = -56'sd1326701376;
localparam signed [55:0] C3_1  = -56'sd1627735824;
localparam signed [55:0] C3_2  =  56'sd3949463232;
localparam signed [55:0] C3_3  =  56'sd1517784840;
localparam signed [55:0] C3_4  = -56'sd3065603112;
localparam signed [55:0] C3_5  = -56'sd461027424;
localparam signed [55:0] C3_6  =  56'sd1234936560;
localparam signed [55:0] C3_7  =  56'sd98583264;
localparam signed [55:0] C3_8  = -56'sd380004768;
localparam signed [55:0] C3_9  = -56'sd13424112;
localparam signed [55:0] C3_10 =  56'sd83779488;
localparam signed [55:0] C3_11 =  56'sd870792;
localparam signed [55:0] C3_12 = -56'sd11694696;
localparam signed [55:0] C3_13 =  56'sd773136;
localparam signed [55:0] C3_14 = -56'sd33700337672601600;

//for c4_scaled
localparam signed [53:0] C4_0  =  54'sd3559107552;
localparam signed [53:0] C4_1  = -54'sd2622761856;
localparam signed [53:0] C4_2  = -54'sd2622761856;
localparam signed [53:0] C4_3  =  54'sd1035288540;
localparam signed [53:0] C4_4  =  54'sd1035288540;
localparam signed [53:0] C4_5  = -54'sd227381440;
localparam signed [53:0] C4_6  = -54'sd227381440;
localparam signed [53:0] C4_7  =  54'sd39721968;
localparam signed [53:0] C4_8  =  54'sd39721968;
localparam signed [53:0] C4_9  = -54'sd4694976;
localparam signed [53:0] C4_10 = -54'sd4694976;
localparam signed [53:0] C4_11 =  54'sd273988;
localparam signed [53:0] C4_12 =  54'sd273988;
localparam signed [53:0] C4_14 = -54'sd4814333953228800;

//for c5_scaled
localparam signed [54:0] C5_0  =  55'sd508443936;
localparam signed [54:0] C5_1  =  55'sd46568808;
localparam signed [54:0] C5_2  = -55'sd936345696;
localparam signed [54:0] C5_3  = -55'sd223836470;
localparam signed [54:0] C5_4  =  55'sd817021062;
localparam signed [54:0] C5_5  =  55'sd121934384;
localparam signed [54:0] C5_6  = -55'sd418526680;
localparam signed [54:0] C5_7  = -55'sd30513912;
localparam signed [54:0] C5_8  =  55'sd138365656;
localparam signed [54:0] C5_9  =  55'sd4453592;
localparam signed [54:0] C5_10 = -55'sd31416528;
localparam signed [54:0] C5_11 = -55'sd300014;
localparam signed [54:0] C5_12 =  55'sd4448158;
localparam signed [54:0] C5_13 = -55'sd296296;
localparam signed [54:0] C5_14 =  55'sd12915289484697600;

//for c6_scaled
localparam signed [51:0] C6_0  = -52'sd534209676;
localparam signed [51:0] C6_1  =  52'sd427901760;
localparam signed [51:0] C6_2  =  52'sd427901760;
localparam signed [51:0] C6_3  = -52'sd217844055;
localparam signed [51:0] C6_4  = -52'sd217844055;
localparam signed [51:0] C6_5  =  52'sd68891680;
localparam signed [51:0] C6_6  =  52'sd68891680;
localparam signed [51:0] C6_7  = -52'sd13406250;
localparam signed [51:0] C6_8  = -52'sd13406250;
localparam signed [51:0] C6_9  =  52'sd1661088;
localparam signed [51:0] C6_10 =  52'sd1661088;
localparam signed [51:0] C6_11 = -52'sd99385;
localparam signed [51:0] C6_12 = -52'sd99385;
localparam signed [51:0] C6_14 =  52'sd1845041354956800;

//for c7_scaled
localparam signed [51:0] C7_0  = -52'sd76315668;
localparam signed [51:0] C7_1  =  52'sd27244503;
localparam signed [51:0] C7_2  =  52'sd106307916;
localparam signed [51:0] C7_3  =  52'sd2371655;
localparam signed [51:0] C7_4  = -52'sd91406601;
localparam signed [51:0] C7_5  = -52'sd6714422;
localparam signed [51:0] C7_6  =  52'sd51231895;
localparam signed [51:0] C7_7  =  52'sd2719002;
localparam signed [51:0] C7_8  = -52'sd18907174;
localparam signed [51:0] C7_9  = -52'sd477191;
localparam signed [51:0] C7_10 =  52'sd4524234;
localparam signed [51:0] C7_11 =  52'sd35321;
localparam signed [51:0] C7_12 = -52'sd657943;
localparam signed [51:0] C7_13 =  52'sd44473;
localparam signed [51:0] C7_14 = -52'sd1938540072268800;

//for c8_scaled
localparam signed [48:0] C8_0  =  49'sd36072036;
localparam signed [48:0] C8_1  = -49'sd29992248;
localparam signed [48:0] C8_2  = -49'sd29992248;
localparam signed [48:0] C8_3  =  49'sd17084925;
localparam signed [48:0] C8_4  =  49'sd17084925;
localparam signed [48:0] C8_5  = -49'sd6477900;
localparam signed [48:0] C8_6  = -49'sd6477900;
localparam signed [48:0] C8_7  =  49'sd1546974;
localparam signed [48:0] C8_8  =  49'sd1546974;
localparam signed [48:0] C8_9  = -49'sd211068;
localparam signed [48:0] C8_10 = -49'sd211068;
localparam signed [48:0] C8_11 =  49'sd13299;
localparam signed [48:0] C8_12 =  49'sd13299;
localparam signed [48:0] C8_14 = -49'sd276934296038400;

//for c9_scaled
localparam signed [47:0] C9_0  =  48'sd5153148;
localparam signed [47:0] C9_1  = -48'sd2938221;
localparam signed [47:0] C9_2  = -48'sd6079788;
localparam signed [47:0] C9_3  =  48'sd1027455;
localparam signed [47:0] C9_4  =  48'sd4984551;
localparam signed [47:0] C9_5  = -48'sd155298;
localparam signed [47:0] C9_6  = -48'sd2850705;
localparam signed [47:0] C9_7  = -48'sd23166;
localparam signed [47:0] C9_8  =  48'sd1116258;
localparam signed [47:0] C9_9  =  48'sd12441;
localparam signed [47:0] C9_10 = -48'sd285714;
localparam signed [47:0] C9_11 = -48'sd1287;
localparam signed [47:0] C9_12 =  48'sd43329;
localparam signed [47:0] C9_13 = -48'sd3003;
localparam signed [47:0] C9_14 =  48'sd130898204236800;

//for c10_scaled
localparam signed [45:0] C10_0  = -46'sd1093092;
localparam signed [45:0] C10_1  =  46'sd926640;
localparam signed [45:0] C10_2  =  46'sd926640;
localparam signed [45:0] C10_3  = -46'sd559845;
localparam signed [45:0] C10_4  = -46'sd559845;
localparam signed [45:0] C10_5  =  46'sd234520;
localparam signed [45:0] C10_6  =  46'sd234520;
localparam signed [45:0] C10_7  = -46'sd64350;
localparam signed [45:0] C10_8  = -46'sd64350;
localparam signed [45:0] C10_9  =  46'sd10296;
localparam signed [45:0] C10_10 =  46'sd10296;
localparam signed [45:0] C10_11 = -46'sd715;
localparam signed [45:0] C10_12 = -46'sd715;
localparam signed [45:0] C10_14 =  46'sd18699743462400;

//for c11_scaled
localparam signed [42:0] C11_0  = -43'sd156156;
localparam signed [42:0] C11_1  =  43'sd106821;
localparam signed [42:0] C11_2  =  43'sd166452;
localparam signed [42:0] C11_3  = -43'sd52195;
localparam signed [42:0] C11_4  = -43'sd129987;
localparam signed [42:0] C11_5  =  43'sd17446;
localparam signed [42:0] C11_6  =  43'sd73645;
localparam signed [42:0] C11_7  = -43'sd3666;
localparam signed [42:0] C11_8  = -43'sd29458;
localparam signed [42:0] C11_9  =  43'sd403;
localparam signed [42:0] C11_10 =  43'sd7878;
localparam signed [42:0] C11_11 = -43'sd13;
localparam signed [42:0] C11_12 = -43'sd1261;
localparam signed [42:0] C11_13 =  43'sd91;
localparam signed [42:0] C11_14 = -43'sd3966612249600;

//for c12_scaled
localparam signed [40:0] C12_0  =  41'sd12012;
localparam signed [40:0] C12_1  = -41'sd10296;
localparam signed [40:0] C12_2  = -41'sd10296;
localparam signed [40:0] C12_3  =  41'sd6435;
localparam signed [40:0] C12_4  =  41'sd6435;
localparam signed [40:0] C12_5  = -41'sd2860;
localparam signed [40:0] C12_6  = -41'sd2860;
localparam signed [40:0] C12_7  =  41'sd858;
localparam signed [40:0] C12_8  =  41'sd858;
localparam signed [40:0] C12_9  = -41'sd156;
localparam signed [40:0] C12_10 = -41'sd156;
localparam signed [40:0] C12_11 =  41'sd13;
localparam signed [40:0] C12_12 =  41'sd13;
localparam signed [40:0] C12_14 = -41'sd566658892800;

//for c13_scaled
localparam signed [36:0] C13_0  =  37'sd1716;
localparam signed [36:0] C13_1  = -37'sd1287;
localparam signed [36:0] C13_2  = -37'sd1716;
localparam signed [36:0] C13_3  =  37'sd715;
localparam signed [36:0] C13_4  =  37'sd1287;
localparam signed [36:0] C13_5  = -37'sd286;
localparam signed [36:0] C13_6  = -37'sd715;
localparam signed [36:0] C13_7  =  37'sd78;
localparam signed [36:0] C13_8  =  37'sd286;
localparam signed [36:0] C13_9  = -37'sd13;
localparam signed [36:0] C13_10 = -37'sd78;
localparam signed [36:0] C13_11 =  37'sd1;
localparam signed [36:0] C13_12 =  37'sd13;
localparam signed [36:0] C13_13 = -37'sd1;
localparam signed [36:0] C13_14 =  37'sd43589145600;
